library verilog;
use verilog.vl_types.all;
entity tstand_vlg_vec_tst is
end tstand_vlg_vec_tst;
