true_S_inst : true_S PORT MAP (
		address	 => address_sig,
		clken	 => clken_sig,
		clock	 => clock_sig,
		q	 => q_sig
	);
