-- ?�N�??N� N�?�???� N??????�N�?�??N� N?N�N�N???N�N?N�?????� ??????N??�?????� ?????�N�?�N�?????????????? N?N?N�N�????N?N�???�
-- N???N?N�??N?N�?�???? ???� N???N�?�???�N?NZN�?�???? ?�??N�?????�N�?� ?????�?? ?? ?????�N�?�N�?????????????? ?�??N�?????�N�?�
-- N???N�?�???�?�?????� ??N?N?N�?�N?N�???�N??�N�N?N? ???� N?N�???????� ??????N�?????????�????


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
library work;
use work.mk_pack.all;			-- ?????????�NZN�?�?�?? ???�???�N�, ?? ????N�??N�???? N??????�N�?�??N�N?N? ???�???�?�N�?�N�??N? N�?????� N????????�?�?� control_y
	
entity Operation_device is					-- ????N�?�N�N�?�??N? ?????�N�?�N�?????????????? N?N?N�N�????N?N�???�
generic(n:integer);			-- ???�N�?�???�N�N� n ?�?�???�?�N� N�?�?�N�N???????N?N�N? N?N?N�N�????N?N�???�
	PORT
	(
		a		:	 IN STD_LOGIC_VECTOR(n-1 DOWNTO 0);	-- 1-N�?? ?????�N�?�???? (???????�???????�)
		b		:	 IN STD_LOGIC_VECTOR(n-1 DOWNTO 0);	-- 2-???? ?????�N�?�???? (???????�??N�?�?�N?)
		clk		:	 IN STD_LOGIC;									--N?????N�N�??N????????�?� 
		set		:	 IN STD_LOGIC;									--N????????�?� ???�N�?�?�N??????? N?N?N�?�??????????
		sno		:	 IN STD_LOGIC;									--N????????�?� ???�N�?�?�?� ?????�N�?�N�????
		sko: out std_logic;											--N????????�?� ??????N�?� ?????�N�?�N�????
		rc		:	 out STD_LOGIC_VECTOR(2*n-1 DOWNTO 0)-- N�?�?�N??�N?N�?�N� (??N�?????�???�???�?????�)
	);
END Operation_device;

architecture behav1 of Operation_device is --??????N??�?????� ?�N�N�??N�?�??N�N????????? N�?�?�?� ?z?? N? ??N??????�N??�?????�?????�?? N?N�N�N???N�N?N�???????? N?N�???�N?
-- ?� ??????N??�?????? ?�N�N�??N�?�??N�N?N�N� ???�???�?�N�??N�N?NZN�N?N? ?????� ?????????????�??N�N� ?z?? ?? ????	

		
component Operation_automat -- ???�???�?�N�?�N�??N? ?????????????�??N�?� ?z??
generic(n:integer);										-- ???�N�?�???�N�N� n ?�?�???�?�N� N�?�?�N�N???????N?N�N? N?N?N�N�????N?N�???�
PORT (y:  in control_y;    								-- N???N�?�???�N?NZN�???� N????????�?�N� ?�?�???�NZN� ??????N�?????????�????N�
	   x: out std_logic_vector(2 downto 0);    		-- ?�??????N�?�N??????� N?N??�??????N?
	   a: in std_logic_vector(n-1 downto 0);    		-- 1-N�?? ?????�N�?�???? (???????�???????�)
	   b: in std_logic_vector(n-1 downto 0);    		-- 2-???? ?????�N�?�???? (???????�??N�?�?�N?)
	   rc: buffer std_logic_vector(2*n-1 downto 0);	-- N�?�?�N??�N?N�?�N� (??N�?????�???�???�?????�)	
	   clk: in std_logic												--N?????N�N�??N????????�?� 
);
end component;

component ControlUnit_meely -- ???�???�?�N�?�N�??N? ?????????????�??N�?� ????
port ( 	
	   y: out control_y;    							--N???N�?�???�N?NZN�???� N????????�?�N�		
	   x: in std_logic_vector(2 downto 0);    	-- ?�??????N�?�N??????� N?N??�??????N?
	   clk: in std_logic;                              --N?????N�N�??N????????�?� 
		set: in std_logic; 										--N????????�?� ???�N�?�?�N??????? N?N?N�?�??????????
		sno: in std_logic;										--N????????�?� ???�N�?�?�?� ?????�N�?�N�????
		sko: out std_logic										--N????????�?� ??????N�?� ?????�N�?�N�????
		);
		end component;
-- ?�?�???�?�N�??N�N??�?? N????????�?�N� ???�N? N????�???????�????N? ?????????????�??N�????		
		
		signal x_X: std_logic_vector(2 downto 0);  		--?�??????N�?�N??????� N?N??�??????N?
		signal y_Y: control_y;									--??????N�?????????�????N�
   
begin	-- ?????�?� ??N�????????N?N�N?N? N????�?�?????�N?N�N� ??????N??�??????, ???�?�??N�?? N????�?�?????�N?N� ?????�?�N� N????????�?�N???N?NZ ???�N�??N?,????N�?�NZN�N?NZ N�???�N? ?�???? ?????�????
unit_OA: Operation_automat				-- unit_OA - N?N�?? ????N? ?z??
GENERIC MAP(n => n
			)					
port map (y_Y,x_X,a,b,rc,clk);		-- ???�N�N�?� ????N�N�???? ???�N? ?z??		
unit_YA: ControlUnit_meely				-- unit_YA - N?N�?? ????N? ????

port map(y=>y_Y,sko=>sko,x=>x_X,clk=>clk,set=>set,sno=>sno);-- ???�N�N�?� ????N�N�???? ???�N? ????

end behav1;