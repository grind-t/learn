library verilog;
use verilog.vl_types.all;
entity Block1_vlg_vec_tst is
end Block1_vlg_vec_tst;
