package mealy_pack is
	type state_s is (s1,s2,s3,s4); 	-- Алфавит состояний
end package mealy_pack;																