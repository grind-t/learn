package pack is							-- Декларация пакета
	type in_x is (x1,x2,x3,x4);      -- Входной алфавит
	type out_y is (y1,y2,y3,y4,y6); 	-- Выходной алфавит
end package pack;							-- Окончание пакета		