library verilog;
use verilog.vl_types.all;
entity automat_myra_vlg_vec_tst is
end automat_myra_vlg_vec_tst;
