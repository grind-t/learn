count_100_inst : count_100 PORT MAP (
		clock	 => clock_sig,
		q	 => q_sig
	);
